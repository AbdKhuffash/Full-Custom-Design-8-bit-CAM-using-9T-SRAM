*** SPICE deck for cell inv{lay} from library CAM8BIT
*** Created on Sat Jul 08, 2023 16:12:20
*** Last revised on Sat Jul 08, 2023 16:17:47
*** Written on Sat Jul 08, 2023 16:17:54 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: inv{lay}
Mnmos@0 out in gnd gnd NMOS L=0.044U W=0.374U AS=0.076P AD=0.063P PS=1.606U PD=1.122U
Mpmos@0 out in vdd vdd PMOS L=0.044U W=0.44U AS=0.086P AD=0.063P PS=1.738U PD=1.122U

* Spice Code nodes in cell cell 'inv{lay}'
vdd vdd 0 DC 1.3
Vin in 0 pulse 1.3 0 0 1p 1p 2n 4n
cload out 0 25fF
.tran 12n
.include D:\rl\22nm.txt
.END
