*** SPICE deck for cell invi{sch} from library invert
*** Created on Fri May 26, 2023 20:31:38
*** Last revised on Fri May 26, 2023 20:35:09
*** Written on Fri May 26, 2023 20:37:30 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT invert__inv FROM CELL inv{sch}
.SUBCKT invert__inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 out in gnd gnd NMOS L=0.4U W=2U
Mpmos@1 vdd in out vdd PMOS L=0.4U W=2U
.ENDS invert__inv

.global gnd vdd

*** TOP LEVEL CELL: invi{sch}
Xinv@0 in out invert__inv

* Spice Code nodes in cell cell 'invi{sch}'
vdd vdd 0 DC 5
vin in 0 pwl 10n 0 20n 5 50n 5 60n 0
cload out 0 250fF
.measure tran tf trig v(out) val=4.5 fall=1 td=8ns trag v(out) val=0.5 fall=1
.measure tran tr trig v(out) val=0.5 rais=1 td=50ns trag v(out) val=4.5 rais=1
.tran 0 0.1us
.include D:\rl\C5_models.txt
.END
