*** SPICE deck for cell nand{lay} from library FullAdder
*** Created on Wed Jun 14, 2023 09:27:55
*** Last revised on Wed Jun 14, 2023 20:47:10
*** Written on Wed Jun 14, 2023 20:47:41 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: nand{lay}
Mnmos@0 gnd a net@47 gnd NMOS L=0.6U W=6U AS=5.4P AD=27P PS=7.8U PD=35.1U
Mnmos@1 net@47 b out gnd NMOS L=0.6U W=6U AS=7.35P AD=5.4P PS=9.5U PD=7.8U
Mpmos@0 vdd a out vdd PMOS L=0.6U W=3U AS=7.35P AD=14.85P PS=9.5U PD=21.3U
Mpmos@1 out b vdd vdd PMOS L=0.6U W=3U AS=14.85P AD=7.35P PS=21.3U PD=9.5U

* Spice Code nodes in cell cell 'nand{lay}'
vdd vdd 0 DC 5
va a 0 pulse 5 0 0 1p 1p 40n 80n
vb b 0 pulse 5 0 0 1p 1p 80n 160n
cload out 0 250fF
.tran 500n
.include D:\rl\C5_models.txt
.END
